package alu_defs;
//--------------------------------------------------------------------
// ALU OPERATIONS
//--------------------------------------------------------------------
	
	parameter ADD =  	3'b000;
	parameter MOV =  	3'b001;
	parameter XOR =   3'b010;
	parameter OR  =  	3'b011;
	parameter SHR =  	3'b100;
	parameter SHL =  	3'b101;
	parameter CMP =   3'b110;
	parameter SUB =   3'b111;
	
endpackage